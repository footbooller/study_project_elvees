package fulladder_env_pkg;

    //uvm_package
    import uvm_pkg::*; 
    import c_pkg::*;
    import fulladder_agent_pkg::*;
    
    `include "uvm_macros.svh"
    `include "fulladder_checker.svh"
    `include "fulladder_env_config.sv"
    `include "fulladder_env.svh"
    //my_package
    
//     `include "fulladder_test.svh"
endpackage:fulladder_env_pkg
