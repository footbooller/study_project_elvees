class fulladder_config extends uvm_object;
    virtual tb_if intf;
endclass