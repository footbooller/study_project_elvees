package fulladder_test_pkg;

    //uvm_package
    import uvm_pkg::*;
    import c_pkg::*;
    import fulladder_agent_pkg::*;
    import fulladder_env_pkg::*;
    
    `include "uvm_macros.svh"
    `include "fulladder_base_test.svh"
    `include "fulladder_test.svh"
    `include "fulladder_cpp_test.svh"
    
endpackage:fulladder_test_pkg
