package fulladder_test_pkg;
    //uvm_package
    import uvm_pkg::*; 
    `include "uvm_macros.svh"
    //my_package
    `include "fulladder_test.svh"
endpackage:fulladder_test_pkg
