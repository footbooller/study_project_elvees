
package c_pkg;
    //uvm_package
    import uvm_pkg::*; 
    `include "uvm_macros.svh"
    //my_package
    `include "base_tr_gen.svh"
endpackage:c_pkg
